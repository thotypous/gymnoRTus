import GetPut::*;
export GetPut::*;
import Clocks::*;
import Reserved::*;
import Connectable::*;
import Vector::*;
import DefaultValue::*;
import MIMO::*;

export DualAD(..);
export DualADWires(..);
export Sample(..);
export ChNum(..);
export ChSample(..);
export mkDualAD;

typedef Bit#(12) Sample;
typedef Bit#(4) ChNum;
typedef Bit#(3) ChSel;
typedef Bit#(8) Byte;

interface DualADWires;
	(* always_ready, result="AD_DIN" *)
	method Bit#(1) getData;
	(* always_ready, enable="AD_SSTRB0", prefix="" *)
	method Action putStrobe0;
	(* always_ready, enable="AD_SSTRB1", prefix="" *)
	method Action putStrobe1;
	(* always_ready, always_enabled, prefix="" *)
	method Action putData0((*port="AD_DOUT0"*)Bit#(1) v);
	(* always_ready, always_enabled, prefix="" *)
	method Action putData1((*port="AD_DOUT1"*)Bit#(1) v);
endinterface

typedef Tuple2#(ChNum, Sample) ChSample;

interface DualAD;
	interface DualADWires wires;
	interface Get#(ChSample) acq;
endinterface

typedef Tuple3#(ChSel, Sample, Sample) InternalTuple;

interface DualADInternal;
	interface DualADWires wires;
	interface Get#(InternalTuple) acq;
endinterface

typedef enum {
	Bipolar  = 1'b0,
	Unipolar = 1'b1
} UniBip deriving (Eq, Bits);

typedef enum {
	Differential = 1'b0,
	SingleEnded  = 1'b1
} SglDif deriving (Eq, Bits);

typedef enum {
	FullPowerDown   = 2'b00,
	FastPowerDown   = 2'b01,
	ReducedPower    = 2'b10,
	NormalOperation = 2'b11
} OperatingMode deriving (Eq, Bits);

// See MAX1280 datasheet p. 14, Table 1
typedef struct {
	ReservedOne#(1) start;
	ChSel sel;
	UniBip unibip;
	SglDif sgldif;
	OperatingMode opmode;
} ControlByte deriving (Eq, Bits);

function Byte makeControlByte(ChSel sel);
	ControlByte ctrl;
	ctrl.sel = sel;
	ctrl.unibip = Unipolar;
	ctrl.sgldif = SingleEnded;
	ctrl.opmode = NormalOperation;
	return pack(ctrl);
endfunction

module mkDualADInternal(DualADInternal);
	// State machine counter
	Array#(Reg#(Bit#(4))) cnt <- mkCReg(3, 0);

	// I/O related
	Reg#(Bit#(1)) din <- mkReg(0);
	Wire#(Bit#(1)) dout0 <- mkWire;
	Wire#(Bit#(1)) dout1 <- mkWire;
	Reg#(Sample) shiftReg0 <- mkRegU;
	Reg#(Sample) shiftReg1 <- mkRegU;

	// Channel and control byte
	Reg#(ChSel) ch <- mkReg(0);
	Reg#(Byte) ctrl <- mkReg(makeControlByte(0));

	// Number of the cycle during which the SSTRB pulse should occur.
	// See MAX1280 datasheet p. 13, Figure 6
	let cycleAfterStrobe = 4'd10;

	// Adjusts the value above considering that there will be an output
	// delay of 2 cycles because of writes to the cnt and din registers.
	let cycleAfterStrobeAdjusted = cycleAfterStrobe + 4'd2;

	(* no_implicit_conditions, fire_when_enabled *)
	rule dinFeed;
		(*split*)
		if (cnt[0] < 8) begin
			// Time to send a bit of the control byte
			din <= ctrl[7];
			ctrl <= ctrl << 1;
		end else begin
			// Time to be quiet
			din <= 0;

			if (cnt[0] == 4'b1111) begin
				// Construct the next control byte
				let nextChannel = ch + 1;
				ctrl <= makeControlByte(nextChannel);
				ch <= nextChannel;
			end
		end
		cnt[0] <= cnt[0] + 1;
	endrule

	let doutBit = cnt[0] - cycleAfterStrobeAdjusted;

	(* fire_when_enabled *)
	rule doutHandle(doutBit < 12);
		shiftReg0 <= (shiftReg0 << 1) | extend(dout0);
		shiftReg1 <= (shiftReg1 << 1) | extend(dout1);
	endrule

	interface DualADWires wires;
		method Bit#(1) getData = din;
		method Action putStrobe0;  cnt[1] <= cycleAfterStrobeAdjusted; endmethod
		method Action putStrobe1;  cnt[2] <= cycleAfterStrobeAdjusted; endmethod
		method Action putData0(v); dout0 <= v; endmethod
		method Action putData1(v); dout1 <= v; endmethod
	endinterface

	interface Get acq;
		method ActionValue#(InternalTuple) get if (doutBit == 12);
			// At the end of the conversion, ch will already be incremented.
			// See MAX1280 datasheet p. 16, Figure 8
			return tuple3(ch - 1, shiftReg0, shiftReg1);
		endmethod
	endinterface
endmodule

module mkDualAD(Clock sClk, DualAD ifc);
	Reset sRst <- mkAsyncResetFromCR(2, sClk);
	let m <- mkDualADInternal(clocked_by sClk, reset_by sRst);

	SyncFIFOIfc#(InternalTuple) sync <- mkSyncFIFOToCC(2, sClk, sRst);
	MIMO#(2, 1, 2, ChSample) mimo <- mkMIMO(defaultValue);

	mkConnection(m.acq, toPut(sync));

	rule mimoPut;
		sync.deq;
		match {.chsel, .sample0, .sample1} = sync.first;
		mimo.enq(2,                           cons(
			tuple2({1'b0, chsel}, sample0),   cons(
			tuple2({1'b1, chsel}, sample1),   nil)
		));
	endrule

	interface wires = m.wires;
	interface Get acq;
		method ActionValue#(ChSample) get;
			mimo.deq(1);
			return mimo.first[0];
		endmethod
	endinterface
endmodule